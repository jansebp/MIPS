module ula(
        input logic [2:0] ULAcontrole,
        input logic a, b,
        input logic cin, addsub, less,
        output logic set, cout,
        output logic ULAsaida
        );

    logic saidaAND, saidaOR, saidaNOR, saidaXOR, saidaADD, saidaSUB, saidaDEF, bAux;
    logic cout0, cout1;

    and ULAand(saidaAND,a,b);                 //000
    or ULAor(saidaOR,a,b);                    //001
    nor ULAnor(saidaNOR,a,b);                 //011
    xor ULAxor(saidaXOR,a,b);                 //101

	 xor ULAaddsub(bAux, b, addsub);
	 adder ULAadd(a, bAux, cin, saidaADD, cout);

    assign set = saidaADD;
	 mux8_1 ULAmux(ULAcontrole, saidaAND, saidaOR, saidaADD, saidaNOR, saidaDEF, saidaXOR, saidaADD, less, ULAsaida);

endmodule
